// Copyright (c) 2017, Yang Zhang, Haipeng Zha, and Huimei Cheng
// All rights reserved.

// Redistribution and use in source and binary forms, with or without
// modification, are permitted provided that the following conditions are met:
    // * Redistributions of source code must retain the above copyright
      // notice, this list of conditions and the following disclaimer.
    // * Redistributions in binary form must reproduce the above copyright
      // notice, this list of conditions and the following disclaimer in the
      // documentation and/or other materials provided with the distribution.
    // * Neither the name of the University of Southern California nor the
      // names of its contributors may be used to endorse or promote products
      // derived from this software without specific prior written permission.

// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL YANG ZHANG, HAIPENG ZHA, AND HUIMEI CHENG BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.




`include "/tools/pdk/stm/.28nm-cmos28fdsoi_24/C28SOI_SC_12_CORE_LR@2.0@20130411.0/behaviour/verilog/C28SOI_SC_12_CORE_LR.v"
`include "/tools/pdk/stm/.28nm-cmos28fdsoi_24/C28SOI_SC_12_CLK_LR@2.1@20130621.0/behaviour/verilog/C28SOI_SC_12_CLK_LR.v"
// In order to run this simulation which includes netlists generated by DC, the above two libraries are supposed to be changed per technology.

 import uvm_pkg::*;
   `include "uvm_macros.svh"
   `include "data_packet.sv"
   `include "edge_driver.sv"
   `include "edge_monitor.sv"
   `include "edge_sequencer.sv"
   `include "edge_agent.sv"
   `include "edge_scoreboard.sv"
   `include "edge_env.sv"
   `include "dut_env.sv"
   `include "edge_sequence_lib.sv"
   `include "test_lib.sv"

module top;   
   bit rst_edge;
   bit rst_edge_ctrl;
   
   bit Lreq;
   bit Rack;
   bit clk;
   wire Lack;
   wire Rreq;

   edge_if ivif(.rst_edge(rst_edge), .rst_edge_ctrl(rst_edge_ctrl), .Rreq(1'b0), .clk(clk));
   edge_if ovif1(.rst_edge(rst_edge), .rst_edge_ctrl(rst_edge_ctrl), .Rreq(1'b0), .clk(clk));
   edge_if ovif2(.rst_edge(rst_edge), .rst_edge_ctrl(rst_edge_ctrl), .Rreq(1'b0), .clk(clk));
   
   // new port: I_SCAN_IN, I_TEST_MODE, I_SCAN_RST, I_SCAN_SE, O_SCAN_OUT
   mlite_cpu_dc uut(.intr_in(ivif.intr_in), .address_next(ovif1.address_next[31:2]), .byte_we_next(ovif1.byte_we_next), .address(ovif1.address[31:2]), .byte_we(ovif1.byte_we), .data_w(ovif1.data_w), .data_r(ivif.data_r), .mem_pause(ivif.mem_pause), .edge_reset(rst_edge), .Lreq(Lreq), .Rack(Rack), .edge_ctrl_reset(rst_edge_ctrl), .Rreq(Rreq), .Lack(Lack), .I_SCAN_IN(1'b0), .I_TEST_MODE(1'b0), .I_SCAN_RST(1'b0), .I_SCAN_SE(1'b0) );
   mlite_cpu_syn uut_ref(.intr_in(ivif.intr_in), .address_next(ovif2.address_next[31:2]), .byte_we_next(ovif2.byte_we_next), .address(ovif2.address[31:2]), .byte_we(ovif2.byte_we), .data_w(ovif2.data_w), .data_r(ivif.data_r), .mem_pause(ivif.mem_pause), .edge_reset(rst_edge), .edge_clk_m(clk), .I_SCAN_IN(1'b0), .I_TEST_MODE(1'b0), .I_SCAN_RST(1'b0), .I_SCAN_SE(1'b0));
   initial begin
      $sdf_annotate("./test/mlite_cpu_dc.sdf",uut,,,"TYPICAL","1.0:1.0:1.0", "FROM_MTM");
      Lreq = 1'b0;
      Rack = 1'b0;
	  clk = 1'b0;

      rst_edge = 1'b1;
      rst_edge_ctrl = 1'b1;
	  
      #5 rst_edge_ctrl = 1'b0;
      #5;
      Lreq = 1'b1;
      wait(Rreq);
      #5 Rack = 1'b1;
	  
      wait(Rreq==0);
      #5 rst_edge_ctrl = 1'b1;
      Lreq = 1'b0;
      Rack = 1'b0;

      #10 rst_edge = 1'b0;
      rst_edge_ctrl = 1'b0;
		
      #50; 
      wait(Rreq != Rack)
      #2;
      Rack = ~Rack;
      forever begin
	Lreq = ~Lreq;
	clk = 1;
	#20; 
	clk = 0;
	wait(Rreq != Rack)
	Rack = ~Rack;
	#20;
      end	
   end

   initial begin
      uvm_config_db#(virtual edge_if)::set(uvm_root::get( ) , "*.agent.*" , "in_intf", ivif);
      uvm_config_db#(virtual edge_if)::set(uvm_root::get( ) , "*.monitor" , "out_intf1", ovif1);
	  uvm_config_db#(virtual edge_if)::set(uvm_root::get( ) , "*.monitor" , "out_intf2", ovif2);
      run_test( );
   end 

endmodule
